entity FRECUENCY_DIVIDER is
PORT (CLK: IN STD_LOGIC;
COUT: OUT STD_LOGIC);
 
end FRECUENCY_DIVIDER;
 
architecture FRECUENCY_DIVIDER_ARCH of FRECUENCY_DIVIDER is
 
SIGNAL Q: STD_LOGIC_VECTOR(23 downto 0);
 
begin
PROCESS(CLK)
BEGIN
IF CLK'EVENT AND CLK = '1' THEN
Q <= Q+1;
END IF;
END PROCESS;
COUT <= Q(17);
end FRECUENCY_DIVIDER_ARCH;
